// Implements a simple Nios II system for the DE-series board.
// Inputs: SW7−0 are parallel port inputs to the Nios II system
// CLOCK_50 is the system clock
// KEY0 is the active-low system reset
// Outputs: LEDR7−0 are parallel port outputs from the Nios II system
module communication (CLOCK_50, SW, KEY, LEDR, dataIn, dataOut);
	input CLOCK_50;
	input [7:0] SW;
	input [0:0] KEY;
	output [9:0] LEDR;

	input dataIn;
	output dataOut;

	assign LEDR[9] = dataIn;
	assign LEDR[8] = dataOut;
	
	wire[31:0] clk;
	clock_divider Divider (CLOCK_50, clk);
	
	wire [7:0] LEDRsub;
	// Instantiate the Nios II system module generated by the Qsys tool:
	nios_system NiosII (
								.charreceived_export(charReceived),    //    charreceived.export
								.charsent_export(charSent),        //        charsent.export
								.clk_clk(CLOCK_50),
								.load_export(load),            //            load.export
								.paralleldatain_export(parallelDataIn),  //  paralleldatain.export
								.paralleldataout_export(parallelDataOut), // paralleldataout.export
								.reset_reset_n(KEY),
								.switches_export(SW),				
								.leds_export(LEDRsub),
								.transen_export(transEn)          //         transen.export
								);
	wire SerialInStart, charReceived, srClockReceive;
	wire [7:0] parallelDataIn;
	
	startBitDetect sbd  (.rst(KEY), .clk(clk[4]), .serialIn(dataIn), .recvStart(SerialInStart), .charRec(charReceived));
	bsc bscRec (.rst(KEY), .clk(clk[4]), .enable(SerialInStart), .srClock(srClockReceive));
	bicReceive bicRec (.rst(KEY), .srClock(srClockReceive), .recEn(SerialInStart), .charRec(charReceived), .clk(clk[4]));
	S2P receiveBuffer (.rst(KEY), .srClock(srClockReceive), .dataIn(dataIn), .data(parallelDataIn));
	
	wire srClockTransmit, transEn, charSent, load;
	wire [7:0] parallelDataOut;
	wire [9:0] p2SBuffer;
	wire [3:0] bitIDCount;
	
	bicTransmit bisTran (.rst(KEY), .srClock(srClockTransmit), .transEn(transEn), .charSent(charSent), .load(load), .clk(clk[4]));
	bsc bscTran (.rst(KEY), .clk(clk[4]), .enable(transEn), .srClock(srClockTransmit));
	P2S transmitBuffer (.rst(KEY), .srClock(srClockTransmit), .data(parallelDataOut), .load(load), .dataOut(dataOut), .transEn(transEn), .clk(clk[4]), .charSent(charSent));
	
	assign LEDR[7:0] = parallelDataIn;
endmodule 
module clock_divider (clock, divided_clocks);
      input   clock;
      output reg [31:0]  divided_clocks;
		
      initial
         divided_clocks = 0;
      always @(posedge clock)
         divided_clocks = divided_clocks + 1;
endmodule
